/* ----------------------------------------------------
 Company : Rochester Institute of Technology (RIT)
 Engineer : Glenn Vodra (GKV4063@rit.edu)

 Create Date : 5/23/23
 Design Name : InstructionMemory
 Module Name : InstructionMemory - dataflow
 Project Name : InstructionFetch

 Description : Mips Instruction Memory
----------------------------------------------------*/

module InstructionMemory(addr, d_out);
	input logic [27:0] addr;
	output logic [31:0] d_out;
	
	//Fibonacci to 10
	logic [7:0] mem [0:371] = '{
		8'h20, 8'h08, 8'h00, 8'h00,
		8'h20, 8'h09, 8'h00, 8'h01,
		8'h20, 8'h0a, 8'h03, 8'hed,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h49, 8'h00, 8'h00,
		8'h01, 8'h28, 8'h40, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h48, 8'h00, 8'h00,
		8'h01, 8'h09, 8'h48, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h49, 8'h00, 8'h00,
		8'h01, 8'h28, 8'h40, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h48, 8'h00, 8'h00,
		8'h01, 8'h09, 8'h48, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h49, 8'h00, 8'h00,
		8'h01, 8'h28, 8'h40, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h48, 8'h00, 8'h00,
		8'h01, 8'h09, 8'h48, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h49, 8'h00, 8'h00,
		8'h01, 8'h28, 8'h40, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h48, 8'h00, 8'h00,
		8'h01, 8'h09, 8'h48, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h49, 8'h00, 8'h00,
		8'h01, 8'h28, 8'h40, 8'h20,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h21, 8'h4a, 8'h00, 8'h01,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'had, 8'h48, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00,
		8'h00, 8'h00, 8'h00, 8'h00
	};
	
	//Acess next four bytes
	always_comb begin
		if (addr < 377) begin
			d_out <= {mem[$unsigned(addr)], mem[$unsigned(addr+1)], mem[$unsigned(addr+2)], mem[$unsigned(addr+3)]};
		end
		else begin
			d_out <= {32{1'b0}};
		end 
	end
	
endmodule
		
