/* ----------------------------------------------------
 Company : Rochester Institute of Technology (RIT)
 Engineer : Glenn Vodra (GKV4063@rit.edu)

 Create Date : 6/5/23

 Package Name : Globals

 Description : Defines N, M and Record Structure 
----------------------------------------------------*/
package global_pkg;
	
	typedef struct {
	//Todo	
	logic a;
	
	}TestRecord;
	
	parameter N = 32;
	parameter M = 5;
	parameter BIT_DEPTH = 32;
	parameter LOG_PORT_DEPTH = 5;
	
endpackage