/* ----------------------------------------------------
 Company : Rochester Institute of Technology (RIT)
 Engineer : Glenn Vodra (GKV4063@rit.edu)

 Create Date : 6/5/23
 Design Name : ExecuteStage
 Module Name : ExecuteStage - Behavioral
 Project Name : RegisterFile

 Description : Execute Stage
----------------------------------------------------*/
//TODO